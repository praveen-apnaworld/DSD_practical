module tb_boolean_exp(
);
reg a,b,c;
wire f1, f2, f3;
boolean_exp uut(a,b,c,f1,f2,f3);
initial begin
a=0; b=0; c=0; #10;
a=0; b=1; c=0; #10;
a=1; b=0; c=1; #10;
a=1; b=1; c=1; #10;
$finish;
end
endmodule

