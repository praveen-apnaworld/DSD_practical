`timescale 1ns / 1ps

module and_gate(
    input a,
    input b,
    output and_gate
);
    assign and_gate = a & b;
endmodule
